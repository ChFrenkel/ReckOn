// Copyright (C) 2020-2022 University of Zurich
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file except in compliance
// with the License, or, at your option, the Apache License version 2.0. You may obtain a copy of the License at
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the License is distributed on
// an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
//------------------------------------------------------------------------------
//
// "lfsr_wout.v" -  Unfolded LFSR module for stochastic updates in output weights
// 
// Project: ReckOn - Spiking RECurrent neural network processor enabling ON-chip learning over second-long timescales
//
// Author:  C. Frenkel, Institute of Neuroinformatics, University of Zurich and ETH Zurich
//
// Cite/paper: [C. Frenkel and G. Indiveri, "ReckOn: A 28nm sub-mm² task-agnostic spiking recurrent neural network
//             processor enabling on-chip learning over second-long timescales," IEEE International Solid-State
//             Circuits Conference (ISSCC), 2022]
//
// Comments: This module has been automatically generated by a custom Python script applying the unfolding algorithm to
//           arbitrary LFSRs (k pseudo-random outputs generated at every clock cycle, where k is the unfolding factor), see 
//               [C. Frenkel, J.D. Legat and D. Bol, "MorphIC: A 65-nm 738k-synapse/mm² quad-core binary-weight digital
//               neuromorphic processor with stochastic spike-driven online learning", IEEE. Trans. on Biomedical Circuits
//               and Systems, vol. 13, no. 5, pp. 999-1010, 2019]
//           for details of the LFSR unfolding procedure.
//
//------------------------------------------------------------------------------


module lfsr_wout (
	// Inputs
	input wire        clk,
	input wire        rst,
	input wire        en,
	input wire [21:0] rst_val,
	input wire [21:0] seed,
	input wire        prog,

	// Output
	output wire [447:0] out
);

	// Nodes definitions
	wire x0, x0a, x0b;
	wire x1, x1a, x1b;
	wire x2, x2a, x2b;
	wire x3, x3a, x3b;
	wire x4, x4a, x4b;
	wire x5, x5a, x5b;
	wire x6, x6a, x6b;
	wire x7, x7a, x7b;
	wire x8, x8a, x8b;
	wire x9, x9a, x9b;
	wire x10, x10a, x10b;
	wire x11, x11a, x11b;
	wire x12, x12a, x12b;
	wire x13, x13a, x13b;
	wire x14, x14a, x14b;
	wire x15, x15a, x15b;
	wire x16, x16a, x16b;
	wire x17, x17a, x17b;
	wire x18, x18a, x18b;
	wire x19, x19a, x19b;
	wire x20, x20a, x20b;
	wire x21, x21a, x21b;
	wire x22, x22a, x22b;
	wire x23, x23a, x23b;
	wire x24, x24a, x24b;
	wire x25, x25a, x25b;
	wire x26, x26a, x26b;
	wire x27, x27a, x27b;
	wire x28, x28a, x28b;
	wire x29, x29a, x29b;
	wire x30, x30a, x30b;
	wire x31, x31a, x31b;
	wire x32, x32a, x32b;
	wire x33, x33a, x33b;
	wire x34, x34a, x34b;
	wire x35, x35a, x35b;
	wire x36, x36a, x36b;
	wire x37, x37a, x37b;
	wire x38, x38a, x38b;
	wire x39, x39a, x39b;
	wire x40, x40a, x40b;
	wire x41, x41a, x41b;
	wire x42, x42a, x42b;
	wire x43, x43a, x43b;
	wire x44, x44a, x44b;
	wire x45, x45a, x45b;
	wire x46, x46a, x46b;
	wire x47, x47a, x47b;
	wire x48, x48a, x48b;
	wire x49, x49a, x49b;
	wire x50, x50a, x50b;
	wire x51, x51a, x51b;
	wire x52, x52a, x52b;
	wire x53, x53a, x53b;
	wire x54, x54a, x54b;
	wire x55, x55a, x55b;
	wire x56, x56a, x56b;
	wire x57, x57a, x57b;
	wire x58, x58a, x58b;
	wire x59, x59a, x59b;
	wire x60, x60a, x60b;
	wire x61, x61a, x61b;
	wire x62, x62a, x62b;
	wire x63, x63a, x63b;
	wire x64, x64a, x64b;
	wire x65, x65a, x65b;
	wire x66, x66a, x66b;
	wire x67, x67a, x67b;
	wire x68, x68a, x68b;
	wire x69, x69a, x69b;
	wire x70, x70a, x70b;
	wire x71, x71a, x71b;
	wire x72, x72a, x72b;
	wire x73, x73a, x73b;
	wire x74, x74a, x74b;
	wire x75, x75a, x75b;
	wire x76, x76a, x76b;
	wire x77, x77a, x77b;
	wire x78, x78a, x78b;
	wire x79, x79a, x79b;
	wire x80, x80a, x80b;
	wire x81, x81a, x81b;
	wire x82, x82a, x82b;
	wire x83, x83a, x83b;
	wire x84, x84a, x84b;
	wire x85, x85a, x85b;
	wire x86, x86a, x86b;
	wire x87, x87a, x87b;
	wire x88, x88a, x88b;
	wire x89, x89a, x89b;
	wire x90, x90a, x90b;
	wire x91, x91a, x91b;
	wire x92, x92a, x92b;
	wire x93, x93a, x93b;
	wire x94, x94a, x94b;
	wire x95, x95a, x95b;
	wire x96, x96a, x96b;
	wire x97, x97a, x97b;
	wire x98, x98a, x98b;
	wire x99, x99a, x99b;
	wire x100, x100a, x100b;
	wire x101, x101a, x101b;
	wire x102, x102a, x102b;
	wire x103, x103a, x103b;
	wire x104, x104a, x104b;
	wire x105, x105a, x105b;
	wire x106, x106a, x106b;
	wire x107, x107a, x107b;
	wire x108, x108a, x108b;
	wire x109, x109a, x109b;
	wire x110, x110a, x110b;
	wire x111, x111a, x111b;
	wire x112, x112a, x112b;
	wire x113, x113a, x113b;
	wire x114, x114a, x114b;
	wire x115, x115a, x115b;
	wire x116, x116a, x116b;
	wire x117, x117a, x117b;
	wire x118, x118a, x118b;
	wire x119, x119a, x119b;
	wire x120, x120a, x120b;
	wire x121, x121a, x121b;
	wire x122, x122a, x122b;
	wire x123, x123a, x123b;
	wire x124, x124a, x124b;
	wire x125, x125a, x125b;
	wire x126, x126a, x126b;
	wire x127, x127a, x127b;
	wire x128, x128a, x128b;
	wire x129, x129a, x129b;
	wire x130, x130a, x130b;
	wire x131, x131a, x131b;
	wire x132, x132a, x132b;
	wire x133, x133a, x133b;
	wire x134, x134a, x134b;
	wire x135, x135a, x135b;
	wire x136, x136a, x136b;
	wire x137, x137a, x137b;
	wire x138, x138a, x138b;
	wire x139, x139a, x139b;
	wire x140, x140a, x140b;
	wire x141, x141a, x141b;
	wire x142, x142a, x142b;
	wire x143, x143a, x143b;
	wire x144, x144a, x144b;
	wire x145, x145a, x145b;
	wire x146, x146a, x146b;
	wire x147, x147a, x147b;
	wire x148, x148a, x148b;
	wire x149, x149a, x149b;
	wire x150, x150a, x150b;
	wire x151, x151a, x151b;
	wire x152, x152a, x152b;
	wire x153, x153a, x153b;
	wire x154, x154a, x154b;
	wire x155, x155a, x155b;
	wire x156, x156a, x156b;
	wire x157, x157a, x157b;
	wire x158, x158a, x158b;
	wire x159, x159a, x159b;
	wire x160, x160a, x160b;
	wire x161, x161a, x161b;
	wire x162, x162a, x162b;
	wire x163, x163a, x163b;
	wire x164, x164a, x164b;
	wire x165, x165a, x165b;
	wire x166, x166a, x166b;
	wire x167, x167a, x167b;
	wire x168, x168a, x168b;
	wire x169, x169a, x169b;
	wire x170, x170a, x170b;
	wire x171, x171a, x171b;
	wire x172, x172a, x172b;
	wire x173, x173a, x173b;
	wire x174, x174a, x174b;
	wire x175, x175a, x175b;
	wire x176, x176a, x176b;
	wire x177, x177a, x177b;
	wire x178, x178a, x178b;
	wire x179, x179a, x179b;
	wire x180, x180a, x180b;
	wire x181, x181a, x181b;
	wire x182, x182a, x182b;
	wire x183, x183a, x183b;
	wire x184, x184a, x184b;
	wire x185, x185a, x185b;
	wire x186, x186a, x186b;
	wire x187, x187a, x187b;
	wire x188, x188a, x188b;
	wire x189, x189a, x189b;
	wire x190, x190a, x190b;
	wire x191, x191a, x191b;
	wire x192, x192a, x192b;
	wire x193, x193a, x193b;
	wire x194, x194a, x194b;
	wire x195, x195a, x195b;
	wire x196, x196a, x196b;
	wire x197, x197a, x197b;
	wire x198, x198a, x198b;
	wire x199, x199a, x199b;
	wire x200, x200a, x200b;
	wire x201, x201a, x201b;
	wire x202, x202a, x202b;
	wire x203, x203a, x203b;
	wire x204, x204a, x204b;
	wire x205, x205a, x205b;
	wire x206, x206a, x206b;
	wire x207, x207a, x207b;
	wire x208, x208a, x208b;
	wire x209, x209a, x209b;
	wire x210, x210a, x210b;
	wire x211, x211a, x211b;
	wire x212, x212a, x212b;
	wire x213, x213a, x213b;
	wire x214, x214a, x214b;
	wire x215, x215a, x215b;
	wire x216, x216a, x216b;
	wire x217, x217a, x217b;
	wire x218, x218a, x218b;
	wire x219, x219a, x219b;
	wire x220, x220a, x220b;
	wire x221, x221a, x221b;
	wire x222, x222a, x222b;
	wire x223, x223a, x223b;
	wire x224, x224a, x224b;
	wire x225, x225a, x225b;
	wire x226, x226a, x226b;
	wire x227, x227a, x227b;
	wire x228, x228a, x228b;
	wire x229, x229a, x229b;
	wire x230, x230a, x230b;
	wire x231, x231a, x231b;
	wire x232, x232a, x232b;
	wire x233, x233a, x233b;
	wire x234, x234a, x234b;
	wire x235, x235a, x235b;
	wire x236, x236a, x236b;
	wire x237, x237a, x237b;
	wire x238, x238a, x238b;
	wire x239, x239a, x239b;
	wire x240, x240a, x240b;
	wire x241, x241a, x241b;
	wire x242, x242a, x242b;
	wire x243, x243a, x243b;
	wire x244, x244a, x244b;
	wire x245, x245a, x245b;
	wire x246, x246a, x246b;
	wire x247, x247a, x247b;
	wire x248, x248a, x248b;
	wire x249, x249a, x249b;
	wire x250, x250a, x250b;
	wire x251, x251a, x251b;
	wire x252, x252a, x252b;
	wire x253, x253a, x253b;
	wire x254, x254a, x254b;
	wire x255, x255a, x255b;
	wire x256, x256a, x256b;
	wire x257, x257a, x257b;
	wire x258, x258a, x258b;
	wire x259, x259a, x259b;
	wire x260, x260a, x260b;
	wire x261, x261a, x261b;
	wire x262, x262a, x262b;
	wire x263, x263a, x263b;
	wire x264, x264a, x264b;
	wire x265, x265a, x265b;
	wire x266, x266a, x266b;
	wire x267, x267a, x267b;
	wire x268, x268a, x268b;
	wire x269, x269a, x269b;
	wire x270, x270a, x270b;
	wire x271, x271a, x271b;
	wire x272, x272a, x272b;
	wire x273, x273a, x273b;
	wire x274, x274a, x274b;
	wire x275, x275a, x275b;
	wire x276, x276a, x276b;
	wire x277, x277a, x277b;
	wire x278, x278a, x278b;
	wire x279, x279a, x279b;
	wire x280, x280a, x280b;
	wire x281, x281a, x281b;
	wire x282, x282a, x282b;
	wire x283, x283a, x283b;
	wire x284, x284a, x284b;
	wire x285, x285a, x285b;
	wire x286, x286a, x286b;
	wire x287, x287a, x287b;
	wire x288, x288a, x288b;
	wire x289, x289a, x289b;
	wire x290, x290a, x290b;
	wire x291, x291a, x291b;
	wire x292, x292a, x292b;
	wire x293, x293a, x293b;
	wire x294, x294a, x294b;
	wire x295, x295a, x295b;
	wire x296, x296a, x296b;
	wire x297, x297a, x297b;
	wire x298, x298a, x298b;
	wire x299, x299a, x299b;
	wire x300, x300a, x300b;
	wire x301, x301a, x301b;
	wire x302, x302a, x302b;
	wire x303, x303a, x303b;
	wire x304, x304a, x304b;
	wire x305, x305a, x305b;
	wire x306, x306a, x306b;
	wire x307, x307a, x307b;
	wire x308, x308a, x308b;
	wire x309, x309a, x309b;
	wire x310, x310a, x310b;
	wire x311, x311a, x311b;
	wire x312, x312a, x312b;
	wire x313, x313a, x313b;
	wire x314, x314a, x314b;
	wire x315, x315a, x315b;
	wire x316, x316a, x316b;
	wire x317, x317a, x317b;
	wire x318, x318a, x318b;
	wire x319, x319a, x319b;
	wire x320, x320a, x320b;
	wire x321, x321a, x321b;
	wire x322, x322a, x322b;
	wire x323, x323a, x323b;
	wire x324, x324a, x324b;
	wire x325, x325a, x325b;
	wire x326, x326a, x326b;
	wire x327, x327a, x327b;
	wire x328, x328a, x328b;
	wire x329, x329a, x329b;
	wire x330, x330a, x330b;
	wire x331, x331a, x331b;
	wire x332, x332a, x332b;
	wire x333, x333a, x333b;
	wire x334, x334a, x334b;
	wire x335, x335a, x335b;
	wire x336, x336a, x336b;
	wire x337, x337a, x337b;
	wire x338, x338a, x338b;
	wire x339, x339a, x339b;
	wire x340, x340a, x340b;
	wire x341, x341a, x341b;
	wire x342, x342a, x342b;
	wire x343, x343a, x343b;
	wire x344, x344a, x344b;
	wire x345, x345a, x345b;
	wire x346, x346a, x346b;
	wire x347, x347a, x347b;
	wire x348, x348a, x348b;
	wire x349, x349a, x349b;
	wire x350, x350a, x350b;
	wire x351, x351a, x351b;
	wire x352, x352a, x352b;
	wire x353, x353a, x353b;
	wire x354, x354a, x354b;
	wire x355, x355a, x355b;
	wire x356, x356a, x356b;
	wire x357, x357a, x357b;
	wire x358, x358a, x358b;
	wire x359, x359a, x359b;
	wire x360, x360a, x360b;
	wire x361, x361a, x361b;
	wire x362, x362a, x362b;
	wire x363, x363a, x363b;
	wire x364, x364a, x364b;
	wire x365, x365a, x365b;
	wire x366, x366a, x366b;
	wire x367, x367a, x367b;
	wire x368, x368a, x368b;
	wire x369, x369a, x369b;
	wire x370, x370a, x370b;
	wire x371, x371a, x371b;
	wire x372, x372a, x372b;
	wire x373, x373a, x373b;
	wire x374, x374a, x374b;
	wire x375, x375a, x375b;
	wire x376, x376a, x376b;
	wire x377, x377a, x377b;
	wire x378, x378a, x378b;
	wire x379, x379a, x379b;
	wire x380, x380a, x380b;
	wire x381, x381a, x381b;
	wire x382, x382a, x382b;
	wire x383, x383a, x383b;
	wire x384, x384a, x384b;
	wire x385, x385a, x385b;
	wire x386, x386a, x386b;
	wire x387, x387a, x387b;
	wire x388, x388a, x388b;
	wire x389, x389a, x389b;
	wire x390, x390a, x390b;
	wire x391, x391a, x391b;
	wire x392, x392a, x392b;
	wire x393, x393a, x393b;
	wire x394, x394a, x394b;
	wire x395, x395a, x395b;
	wire x396, x396a, x396b;
	wire x397, x397a, x397b;
	wire x398, x398a, x398b;
	wire x399, x399a, x399b;
	wire x400, x400a, x400b;
	wire x401, x401a, x401b;
	wire x402, x402a, x402b;
	wire x403, x403a, x403b;
	wire x404, x404a, x404b;
	wire x405, x405a, x405b;
	wire x406, x406a, x406b;
	wire x407, x407a, x407b;
	wire x408, x408a, x408b;
	wire x409, x409a, x409b;
	wire x410, x410a, x410b;
	wire x411, x411a, x411b;
	wire x412, x412a, x412b;
	wire x413, x413a, x413b;
	wire x414, x414a, x414b;
	wire x415, x415a, x415b;
	wire x416, x416a, x416b;
	wire x417, x417a, x417b;
	wire x418, x418a, x418b;
	wire x419, x419a, x419b;
	wire x420, x420a, x420b;
	wire x421, x421a, x421b;
	wire x422, x422a, x422b;
	wire x423, x423a, x423b;
	wire x424, x424a, x424b;
	wire x425, x425a, x425b;
	wire x426, x426a, x426b;
	wire x427, x427a, x427b;
	wire x428, x428a, x428b;
	wire x429, x429a, x429b;
	wire x430, x430a, x430b;
	wire x431, x431a, x431b;
	wire x432, x432a, x432b;
	wire x433, x433a, x433b;
	wire x434, x434a, x434b;
	wire x435, x435a, x435b;
	wire x436, x436a, x436b;
	wire x437, x437a, x437b;
	wire x438, x438a, x438b;
	wire x439, x439a, x439b;
	wire x440, x440a, x440b;
	wire x441, x441a, x441b;
	wire x442, x442a, x442b;
	wire x443, x443a, x443b;
	wire x444, x444a, x444b;
	wire x445, x445a, x445b;
	wire x446, x446a, x446b;
	wire x447, x447a, x447b;
	wire y0;
	wire y1;
	wire y2;
	wire y3;
	wire y4;
	wire y5;
	wire y6;
	wire y7;
	wire y8;
	wire y9;
	wire y10;
	wire y11;
	wire y12;
	wire y13;
	wire y14;
	wire y15;
	wire y16;
	wire y17;
	wire y18;
	wire y19;
	wire y20;
	wire y21;
	wire y22;
	wire y23;
	wire y24;
	wire y25;
	wire y26;
	wire y27;
	wire y28;
	wire y29;
	wire y30;
	wire y31;
	wire y32;
	wire y33;
	wire y34;
	wire y35;
	wire y36;
	wire y37;
	wire y38;
	wire y39;
	wire y40;
	wire y41;
	wire y42;
	wire y43;
	wire y44;
	wire y45;
	wire y46;
	wire y47;
	wire y48;
	wire y49;
	wire y50;
	wire y51;
	wire y52;
	wire y53;
	wire y54;
	wire y55;
	wire y56;
	wire y57;
	wire y58;
	wire y59;
	wire y60;
	wire y61;
	wire y62;
	wire y63;
	wire y64;
	wire y65;
	wire y66;
	wire y67;
	wire y68;
	wire y69;
	wire y70;
	wire y71;
	wire y72;
	wire y73;
	wire y74;
	wire y75;
	wire y76;
	wire y77;
	wire y78;
	wire y79;
	wire y80;
	wire y81;
	wire y82;
	wire y83;
	wire y84;
	wire y85;
	wire y86;
	wire y87;
	wire y88;
	wire y89;
	wire y90;
	wire y91;
	wire y92;
	wire y93;
	wire y94;
	wire y95;
	wire y96;
	wire y97;
	wire y98;
	wire y99;
	wire y100;
	wire y101;
	wire y102;
	wire y103;
	wire y104;
	wire y105;
	wire y106;
	wire y107;
	wire y108;
	wire y109;
	wire y110;
	wire y111;
	wire y112;
	wire y113;
	wire y114;
	wire y115;
	wire y116;
	wire y117;
	wire y118;
	wire y119;
	wire y120;
	wire y121;
	wire y122;
	wire y123;
	wire y124;
	wire y125;
	wire y126;
	wire y127;
	wire y128;
	wire y129;
	wire y130;
	wire y131;
	wire y132;
	wire y133;
	wire y134;
	wire y135;
	wire y136;
	wire y137;
	wire y138;
	wire y139;
	wire y140;
	wire y141;
	wire y142;
	wire y143;
	wire y144;
	wire y145;
	wire y146;
	wire y147;
	wire y148;
	wire y149;
	wire y150;
	wire y151;
	wire y152;
	wire y153;
	wire y154;
	wire y155;
	wire y156;
	wire y157;
	wire y158;
	wire y159;
	wire y160;
	wire y161;
	wire y162;
	wire y163;
	wire y164;
	wire y165;
	wire y166;
	wire y167;
	wire y168;
	wire y169;
	wire y170;
	wire y171;
	wire y172;
	wire y173;
	wire y174;
	wire y175;
	wire y176;
	wire y177;
	wire y178;
	wire y179;
	wire y180;
	wire y181;
	wire y182;
	wire y183;
	wire y184;
	wire y185;
	wire y186;
	wire y187;
	wire y188;
	wire y189;
	wire y190;
	wire y191;
	wire y192;
	wire y193;
	wire y194;
	wire y195;
	wire y196;
	wire y197;
	wire y198;
	wire y199;
	wire y200;
	wire y201;
	wire y202;
	wire y203;
	wire y204;
	wire y205;
	wire y206;
	wire y207;
	wire y208;
	wire y209;
	wire y210;
	wire y211;
	wire y212;
	wire y213;
	wire y214;
	wire y215;
	wire y216;
	wire y217;
	wire y218;
	wire y219;
	wire y220;
	wire y221;
	wire y222;
	wire y223;
	wire y224;
	wire y225;
	wire y226;
	wire y227;
	wire y228;
	wire y229;
	wire y230;
	wire y231;
	wire y232;
	wire y233;
	wire y234;
	wire y235;
	wire y236;
	wire y237;
	wire y238;
	wire y239;
	wire y240;
	wire y241;
	wire y242;
	wire y243;
	wire y244;
	wire y245;
	wire y246;
	wire y247;
	wire y248;
	wire y249;
	wire y250;
	wire y251;
	wire y252;
	wire y253;
	wire y254;
	wire y255;
	wire y256;
	wire y257;
	wire y258;
	wire y259;
	wire y260;
	wire y261;
	wire y262;
	wire y263;
	wire y264;
	wire y265;
	wire y266;
	wire y267;
	wire y268;
	wire y269;
	wire y270;
	wire y271;
	wire y272;
	wire y273;
	wire y274;
	wire y275;
	wire y276;
	wire y277;
	wire y278;
	wire y279;
	wire y280;
	wire y281;
	wire y282;
	wire y283;
	wire y284;
	wire y285;
	wire y286;
	wire y287;
	wire y288;
	wire y289;
	wire y290;
	wire y291;
	wire y292;
	wire y293;
	wire y294;
	wire y295;
	wire y296;
	wire y297;
	wire y298;
	wire y299;
	wire y300;
	wire y301;
	wire y302;
	wire y303;
	wire y304;
	wire y305;
	wire y306;
	wire y307;
	wire y308;
	wire y309;
	wire y310;
	wire y311;
	wire y312;
	wire y313;
	wire y314;
	wire y315;
	wire y316;
	wire y317;
	wire y318;
	wire y319;
	wire y320;
	wire y321;
	wire y322;
	wire y323;
	wire y324;
	wire y325;
	wire y326;
	wire y327;
	wire y328;
	wire y329;
	wire y330;
	wire y331;
	wire y332;
	wire y333;
	wire y334;
	wire y335;
	wire y336;
	wire y337;
	wire y338;
	wire y339;
	wire y340;
	wire y341;
	wire y342;
	wire y343;
	wire y344;
	wire y345;
	wire y346;
	wire y347;
	wire y348;
	wire y349;
	wire y350;
	wire y351;
	wire y352;
	wire y353;
	wire y354;
	wire y355;
	wire y356;
	wire y357;
	wire y358;
	wire y359;
	wire y360;
	wire y361;
	wire y362;
	wire y363;
	wire y364;
	wire y365;
	wire y366;
	wire y367;
	wire y368;
	wire y369;
	wire y370;
	wire y371;
	wire y372;
	wire y373;
	wire y374;
	wire y375;
	wire y376;
	wire y377;
	wire y378;
	wire y379;
	wire y380;
	wire y381;
	wire y382;
	wire y383;
	wire y384;
	wire y385;
	wire y386;
	wire y387;
	wire y388;
	wire y389;
	wire y390;
	wire y391;
	wire y392;
	wire y393;
	wire y394;
	wire y395;
	wire y396;
	wire y397;
	wire y398;
	wire y399;
	wire y400;
	wire y401;
	wire y402;
	wire y403;
	wire y404;
	wire y405;
	wire y406;
	wire y407;
	wire y408;
	wire y409;
	wire y410;
	wire y411;
	wire y412;
	wire y413;
	wire y414;
	wire y415;
	wire y416;
	wire y417;
	wire y418;
	wire y419;
	wire y420;
	wire y421;
	wire y422;
	wire y423;
	wire y424;
	wire y425;
	wire y426;
	wire y427;
	wire y428;
	wire y429;
	wire y430;
	wire y431;
	wire y432;
	wire y433;
	wire y434;
	wire y435;
	wire y436;
	wire y437;
	wire y438;
	wire y439;
	wire y440;
	wire y441;
	wire y442;
	wire y443;
	wire y444;
	wire y445;
	wire y446;
	wire y447;
	reg d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21;

	// Combinational and sequential logic definitions
	assign x0 = x0a ^ x0b;
	assign x1 = x1a ^ x1b;
	assign x2 = x2a ^ x2b;
	assign x3 = x3a ^ x3b;
	assign x4 = x4a ^ x4b;
	assign x5 = x5a ^ x5b;
	assign x6 = x6a ^ x6b;
	assign x7 = x7a ^ x7b;
	assign x8 = x8a ^ x8b;
	assign x9 = x9a ^ x9b;
	assign x10 = x10a ^ x10b;
	assign x11 = x11a ^ x11b;
	assign x12 = x12a ^ x12b;
	assign x13 = x13a ^ x13b;
	assign x14 = x14a ^ x14b;
	assign x15 = x15a ^ x15b;
	assign x16 = x16a ^ x16b;
	assign x17 = x17a ^ x17b;
	assign x18 = x18a ^ x18b;
	assign x19 = x19a ^ x19b;
	assign x20 = x20a ^ x20b;
	assign x21 = x21a ^ x21b;
	assign x22 = x22a ^ x22b;
	assign x23 = x23a ^ x23b;
	assign x24 = x24a ^ x24b;
	assign x25 = x25a ^ x25b;
	assign x26 = x26a ^ x26b;
	assign x27 = x27a ^ x27b;
	assign x28 = x28a ^ x28b;
	assign x29 = x29a ^ x29b;
	assign x30 = x30a ^ x30b;
	assign x31 = x31a ^ x31b;
	assign x32 = x32a ^ x32b;
	assign x33 = x33a ^ x33b;
	assign x34 = x34a ^ x34b;
	assign x35 = x35a ^ x35b;
	assign x36 = x36a ^ x36b;
	assign x37 = x37a ^ x37b;
	assign x38 = x38a ^ x38b;
	assign x39 = x39a ^ x39b;
	assign x40 = x40a ^ x40b;
	assign x41 = x41a ^ x41b;
	assign x42 = x42a ^ x42b;
	assign x43 = x43a ^ x43b;
	assign x44 = x44a ^ x44b;
	assign x45 = x45a ^ x45b;
	assign x46 = x46a ^ x46b;
	assign x47 = x47a ^ x47b;
	assign x48 = x48a ^ x48b;
	assign x49 = x49a ^ x49b;
	assign x50 = x50a ^ x50b;
	assign x51 = x51a ^ x51b;
	assign x52 = x52a ^ x52b;
	assign x53 = x53a ^ x53b;
	assign x54 = x54a ^ x54b;
	assign x55 = x55a ^ x55b;
	assign x56 = x56a ^ x56b;
	assign x57 = x57a ^ x57b;
	assign x58 = x58a ^ x58b;
	assign x59 = x59a ^ x59b;
	assign x60 = x60a ^ x60b;
	assign x61 = x61a ^ x61b;
	assign x62 = x62a ^ x62b;
	assign x63 = x63a ^ x63b;
	assign x64 = x64a ^ x64b;
	assign x65 = x65a ^ x65b;
	assign x66 = x66a ^ x66b;
	assign x67 = x67a ^ x67b;
	assign x68 = x68a ^ x68b;
	assign x69 = x69a ^ x69b;
	assign x70 = x70a ^ x70b;
	assign x71 = x71a ^ x71b;
	assign x72 = x72a ^ x72b;
	assign x73 = x73a ^ x73b;
	assign x74 = x74a ^ x74b;
	assign x75 = x75a ^ x75b;
	assign x76 = x76a ^ x76b;
	assign x77 = x77a ^ x77b;
	assign x78 = x78a ^ x78b;
	assign x79 = x79a ^ x79b;
	assign x80 = x80a ^ x80b;
	assign x81 = x81a ^ x81b;
	assign x82 = x82a ^ x82b;
	assign x83 = x83a ^ x83b;
	assign x84 = x84a ^ x84b;
	assign x85 = x85a ^ x85b;
	assign x86 = x86a ^ x86b;
	assign x87 = x87a ^ x87b;
	assign x88 = x88a ^ x88b;
	assign x89 = x89a ^ x89b;
	assign x90 = x90a ^ x90b;
	assign x91 = x91a ^ x91b;
	assign x92 = x92a ^ x92b;
	assign x93 = x93a ^ x93b;
	assign x94 = x94a ^ x94b;
	assign x95 = x95a ^ x95b;
	assign x96 = x96a ^ x96b;
	assign x97 = x97a ^ x97b;
	assign x98 = x98a ^ x98b;
	assign x99 = x99a ^ x99b;
	assign x100 = x100a ^ x100b;
	assign x101 = x101a ^ x101b;
	assign x102 = x102a ^ x102b;
	assign x103 = x103a ^ x103b;
	assign x104 = x104a ^ x104b;
	assign x105 = x105a ^ x105b;
	assign x106 = x106a ^ x106b;
	assign x107 = x107a ^ x107b;
	assign x108 = x108a ^ x108b;
	assign x109 = x109a ^ x109b;
	assign x110 = x110a ^ x110b;
	assign x111 = x111a ^ x111b;
	assign x112 = x112a ^ x112b;
	assign x113 = x113a ^ x113b;
	assign x114 = x114a ^ x114b;
	assign x115 = x115a ^ x115b;
	assign x116 = x116a ^ x116b;
	assign x117 = x117a ^ x117b;
	assign x118 = x118a ^ x118b;
	assign x119 = x119a ^ x119b;
	assign x120 = x120a ^ x120b;
	assign x121 = x121a ^ x121b;
	assign x122 = x122a ^ x122b;
	assign x123 = x123a ^ x123b;
	assign x124 = x124a ^ x124b;
	assign x125 = x125a ^ x125b;
	assign x126 = x126a ^ x126b;
	assign x127 = x127a ^ x127b;
	assign x128 = x128a ^ x128b;
	assign x129 = x129a ^ x129b;
	assign x130 = x130a ^ x130b;
	assign x131 = x131a ^ x131b;
	assign x132 = x132a ^ x132b;
	assign x133 = x133a ^ x133b;
	assign x134 = x134a ^ x134b;
	assign x135 = x135a ^ x135b;
	assign x136 = x136a ^ x136b;
	assign x137 = x137a ^ x137b;
	assign x138 = x138a ^ x138b;
	assign x139 = x139a ^ x139b;
	assign x140 = x140a ^ x140b;
	assign x141 = x141a ^ x141b;
	assign x142 = x142a ^ x142b;
	assign x143 = x143a ^ x143b;
	assign x144 = x144a ^ x144b;
	assign x145 = x145a ^ x145b;
	assign x146 = x146a ^ x146b;
	assign x147 = x147a ^ x147b;
	assign x148 = x148a ^ x148b;
	assign x149 = x149a ^ x149b;
	assign x150 = x150a ^ x150b;
	assign x151 = x151a ^ x151b;
	assign x152 = x152a ^ x152b;
	assign x153 = x153a ^ x153b;
	assign x154 = x154a ^ x154b;
	assign x155 = x155a ^ x155b;
	assign x156 = x156a ^ x156b;
	assign x157 = x157a ^ x157b;
	assign x158 = x158a ^ x158b;
	assign x159 = x159a ^ x159b;
	assign x160 = x160a ^ x160b;
	assign x161 = x161a ^ x161b;
	assign x162 = x162a ^ x162b;
	assign x163 = x163a ^ x163b;
	assign x164 = x164a ^ x164b;
	assign x165 = x165a ^ x165b;
	assign x166 = x166a ^ x166b;
	assign x167 = x167a ^ x167b;
	assign x168 = x168a ^ x168b;
	assign x169 = x169a ^ x169b;
	assign x170 = x170a ^ x170b;
	assign x171 = x171a ^ x171b;
	assign x172 = x172a ^ x172b;
	assign x173 = x173a ^ x173b;
	assign x174 = x174a ^ x174b;
	assign x175 = x175a ^ x175b;
	assign x176 = x176a ^ x176b;
	assign x177 = x177a ^ x177b;
	assign x178 = x178a ^ x178b;
	assign x179 = x179a ^ x179b;
	assign x180 = x180a ^ x180b;
	assign x181 = x181a ^ x181b;
	assign x182 = x182a ^ x182b;
	assign x183 = x183a ^ x183b;
	assign x184 = x184a ^ x184b;
	assign x185 = x185a ^ x185b;
	assign x186 = x186a ^ x186b;
	assign x187 = x187a ^ x187b;
	assign x188 = x188a ^ x188b;
	assign x189 = x189a ^ x189b;
	assign x190 = x190a ^ x190b;
	assign x191 = x191a ^ x191b;
	assign x192 = x192a ^ x192b;
	assign x193 = x193a ^ x193b;
	assign x194 = x194a ^ x194b;
	assign x195 = x195a ^ x195b;
	assign x196 = x196a ^ x196b;
	assign x197 = x197a ^ x197b;
	assign x198 = x198a ^ x198b;
	assign x199 = x199a ^ x199b;
	assign x200 = x200a ^ x200b;
	assign x201 = x201a ^ x201b;
	assign x202 = x202a ^ x202b;
	assign x203 = x203a ^ x203b;
	assign x204 = x204a ^ x204b;
	assign x205 = x205a ^ x205b;
	assign x206 = x206a ^ x206b;
	assign x207 = x207a ^ x207b;
	assign x208 = x208a ^ x208b;
	assign x209 = x209a ^ x209b;
	assign x210 = x210a ^ x210b;
	assign x211 = x211a ^ x211b;
	assign x212 = x212a ^ x212b;
	assign x213 = x213a ^ x213b;
	assign x214 = x214a ^ x214b;
	assign x215 = x215a ^ x215b;
	assign x216 = x216a ^ x216b;
	assign x217 = x217a ^ x217b;
	assign x218 = x218a ^ x218b;
	assign x219 = x219a ^ x219b;
	assign x220 = x220a ^ x220b;
	assign x221 = x221a ^ x221b;
	assign x222 = x222a ^ x222b;
	assign x223 = x223a ^ x223b;
	assign x224 = x224a ^ x224b;
	assign x225 = x225a ^ x225b;
	assign x226 = x226a ^ x226b;
	assign x227 = x227a ^ x227b;
	assign x228 = x228a ^ x228b;
	assign x229 = x229a ^ x229b;
	assign x230 = x230a ^ x230b;
	assign x231 = x231a ^ x231b;
	assign x232 = x232a ^ x232b;
	assign x233 = x233a ^ x233b;
	assign x234 = x234a ^ x234b;
	assign x235 = x235a ^ x235b;
	assign x236 = x236a ^ x236b;
	assign x237 = x237a ^ x237b;
	assign x238 = x238a ^ x238b;
	assign x239 = x239a ^ x239b;
	assign x240 = x240a ^ x240b;
	assign x241 = x241a ^ x241b;
	assign x242 = x242a ^ x242b;
	assign x243 = x243a ^ x243b;
	assign x244 = x244a ^ x244b;
	assign x245 = x245a ^ x245b;
	assign x246 = x246a ^ x246b;
	assign x247 = x247a ^ x247b;
	assign x248 = x248a ^ x248b;
	assign x249 = x249a ^ x249b;
	assign x250 = x250a ^ x250b;
	assign x251 = x251a ^ x251b;
	assign x252 = x252a ^ x252b;
	assign x253 = x253a ^ x253b;
	assign x254 = x254a ^ x254b;
	assign x255 = x255a ^ x255b;
	assign x256 = x256a ^ x256b;
	assign x257 = x257a ^ x257b;
	assign x258 = x258a ^ x258b;
	assign x259 = x259a ^ x259b;
	assign x260 = x260a ^ x260b;
	assign x261 = x261a ^ x261b;
	assign x262 = x262a ^ x262b;
	assign x263 = x263a ^ x263b;
	assign x264 = x264a ^ x264b;
	assign x265 = x265a ^ x265b;
	assign x266 = x266a ^ x266b;
	assign x267 = x267a ^ x267b;
	assign x268 = x268a ^ x268b;
	assign x269 = x269a ^ x269b;
	assign x270 = x270a ^ x270b;
	assign x271 = x271a ^ x271b;
	assign x272 = x272a ^ x272b;
	assign x273 = x273a ^ x273b;
	assign x274 = x274a ^ x274b;
	assign x275 = x275a ^ x275b;
	assign x276 = x276a ^ x276b;
	assign x277 = x277a ^ x277b;
	assign x278 = x278a ^ x278b;
	assign x279 = x279a ^ x279b;
	assign x280 = x280a ^ x280b;
	assign x281 = x281a ^ x281b;
	assign x282 = x282a ^ x282b;
	assign x283 = x283a ^ x283b;
	assign x284 = x284a ^ x284b;
	assign x285 = x285a ^ x285b;
	assign x286 = x286a ^ x286b;
	assign x287 = x287a ^ x287b;
	assign x288 = x288a ^ x288b;
	assign x289 = x289a ^ x289b;
	assign x290 = x290a ^ x290b;
	assign x291 = x291a ^ x291b;
	assign x292 = x292a ^ x292b;
	assign x293 = x293a ^ x293b;
	assign x294 = x294a ^ x294b;
	assign x295 = x295a ^ x295b;
	assign x296 = x296a ^ x296b;
	assign x297 = x297a ^ x297b;
	assign x298 = x298a ^ x298b;
	assign x299 = x299a ^ x299b;
	assign x300 = x300a ^ x300b;
	assign x301 = x301a ^ x301b;
	assign x302 = x302a ^ x302b;
	assign x303 = x303a ^ x303b;
	assign x304 = x304a ^ x304b;
	assign x305 = x305a ^ x305b;
	assign x306 = x306a ^ x306b;
	assign x307 = x307a ^ x307b;
	assign x308 = x308a ^ x308b;
	assign x309 = x309a ^ x309b;
	assign x310 = x310a ^ x310b;
	assign x311 = x311a ^ x311b;
	assign x312 = x312a ^ x312b;
	assign x313 = x313a ^ x313b;
	assign x314 = x314a ^ x314b;
	assign x315 = x315a ^ x315b;
	assign x316 = x316a ^ x316b;
	assign x317 = x317a ^ x317b;
	assign x318 = x318a ^ x318b;
	assign x319 = x319a ^ x319b;
	assign x320 = x320a ^ x320b;
	assign x321 = x321a ^ x321b;
	assign x322 = x322a ^ x322b;
	assign x323 = x323a ^ x323b;
	assign x324 = x324a ^ x324b;
	assign x325 = x325a ^ x325b;
	assign x326 = x326a ^ x326b;
	assign x327 = x327a ^ x327b;
	assign x328 = x328a ^ x328b;
	assign x329 = x329a ^ x329b;
	assign x330 = x330a ^ x330b;
	assign x331 = x331a ^ x331b;
	assign x332 = x332a ^ x332b;
	assign x333 = x333a ^ x333b;
	assign x334 = x334a ^ x334b;
	assign x335 = x335a ^ x335b;
	assign x336 = x336a ^ x336b;
	assign x337 = x337a ^ x337b;
	assign x338 = x338a ^ x338b;
	assign x339 = x339a ^ x339b;
	assign x340 = x340a ^ x340b;
	assign x341 = x341a ^ x341b;
	assign x342 = x342a ^ x342b;
	assign x343 = x343a ^ x343b;
	assign x344 = x344a ^ x344b;
	assign x345 = x345a ^ x345b;
	assign x346 = x346a ^ x346b;
	assign x347 = x347a ^ x347b;
	assign x348 = x348a ^ x348b;
	assign x349 = x349a ^ x349b;
	assign x350 = x350a ^ x350b;
	assign x351 = x351a ^ x351b;
	assign x352 = x352a ^ x352b;
	assign x353 = x353a ^ x353b;
	assign x354 = x354a ^ x354b;
	assign x355 = x355a ^ x355b;
	assign x356 = x356a ^ x356b;
	assign x357 = x357a ^ x357b;
	assign x358 = x358a ^ x358b;
	assign x359 = x359a ^ x359b;
	assign x360 = x360a ^ x360b;
	assign x361 = x361a ^ x361b;
	assign x362 = x362a ^ x362b;
	assign x363 = x363a ^ x363b;
	assign x364 = x364a ^ x364b;
	assign x365 = x365a ^ x365b;
	assign x366 = x366a ^ x366b;
	assign x367 = x367a ^ x367b;
	assign x368 = x368a ^ x368b;
	assign x369 = x369a ^ x369b;
	assign x370 = x370a ^ x370b;
	assign x371 = x371a ^ x371b;
	assign x372 = x372a ^ x372b;
	assign x373 = x373a ^ x373b;
	assign x374 = x374a ^ x374b;
	assign x375 = x375a ^ x375b;
	assign x376 = x376a ^ x376b;
	assign x377 = x377a ^ x377b;
	assign x378 = x378a ^ x378b;
	assign x379 = x379a ^ x379b;
	assign x380 = x380a ^ x380b;
	assign x381 = x381a ^ x381b;
	assign x382 = x382a ^ x382b;
	assign x383 = x383a ^ x383b;
	assign x384 = x384a ^ x384b;
	assign x385 = x385a ^ x385b;
	assign x386 = x386a ^ x386b;
	assign x387 = x387a ^ x387b;
	assign x388 = x388a ^ x388b;
	assign x389 = x389a ^ x389b;
	assign x390 = x390a ^ x390b;
	assign x391 = x391a ^ x391b;
	assign x392 = x392a ^ x392b;
	assign x393 = x393a ^ x393b;
	assign x394 = x394a ^ x394b;
	assign x395 = x395a ^ x395b;
	assign x396 = x396a ^ x396b;
	assign x397 = x397a ^ x397b;
	assign x398 = x398a ^ x398b;
	assign x399 = x399a ^ x399b;
	assign x400 = x400a ^ x400b;
	assign x401 = x401a ^ x401b;
	assign x402 = x402a ^ x402b;
	assign x403 = x403a ^ x403b;
	assign x404 = x404a ^ x404b;
	assign x405 = x405a ^ x405b;
	assign x406 = x406a ^ x406b;
	assign x407 = x407a ^ x407b;
	assign x408 = x408a ^ x408b;
	assign x409 = x409a ^ x409b;
	assign x410 = x410a ^ x410b;
	assign x411 = x411a ^ x411b;
	assign x412 = x412a ^ x412b;
	assign x413 = x413a ^ x413b;
	assign x414 = x414a ^ x414b;
	assign x415 = x415a ^ x415b;
	assign x416 = x416a ^ x416b;
	assign x417 = x417a ^ x417b;
	assign x418 = x418a ^ x418b;
	assign x419 = x419a ^ x419b;
	assign x420 = x420a ^ x420b;
	assign x421 = x421a ^ x421b;
	assign x422 = x422a ^ x422b;
	assign x423 = x423a ^ x423b;
	assign x424 = x424a ^ x424b;
	assign x425 = x425a ^ x425b;
	assign x426 = x426a ^ x426b;
	assign x427 = x427a ^ x427b;
	assign x428 = x428a ^ x428b;
	assign x429 = x429a ^ x429b;
	assign x430 = x430a ^ x430b;
	assign x431 = x431a ^ x431b;
	assign x432 = x432a ^ x432b;
	assign x433 = x433a ^ x433b;
	assign x434 = x434a ^ x434b;
	assign x435 = x435a ^ x435b;
	assign x436 = x436a ^ x436b;
	assign x437 = x437a ^ x437b;
	assign x438 = x438a ^ x438b;
	assign x439 = x439a ^ x439b;
	assign x440 = x440a ^ x440b;
	assign x441 = x441a ^ x441b;
	assign x442 = x442a ^ x442b;
	assign x443 = x443a ^ x443b;
	assign x444 = x444a ^ x444b;
	assign x445 = x445a ^ x445b;
	assign x446 = x446a ^ x446b;
	assign x447 = x447a ^ x447b;
	assign y1 = x0;
	assign y2 = x1;
	assign y3 = x2;
	assign y4 = x3;
	assign y5 = x4;
	assign y6 = x5;
	assign y7 = x6;
	assign y8 = x7;
	assign y9 = x8;
	assign y10 = x9;
	assign y11 = x10;
	assign y12 = x11;
	assign y13 = x12;
	assign y14 = x13;
	assign y15 = x14;
	assign y16 = x15;
	assign y17 = x16;
	assign y18 = x17;
	assign y19 = x18;
	assign y20 = x19;
	assign y21 = x20;
	assign y22 = x21;
	assign y23 = x22;
	assign y24 = x23;
	assign y25 = x24;
	assign y26 = x25;
	assign y27 = x26;
	assign y28 = x27;
	assign y29 = x28;
	assign y30 = x29;
	assign y31 = x30;
	assign y32 = x31;
	assign y33 = x32;
	assign y34 = x33;
	assign y35 = x34;
	assign y36 = x35;
	assign y37 = x36;
	assign y38 = x37;
	assign y39 = x38;
	assign y40 = x39;
	assign y41 = x40;
	assign y42 = x41;
	assign y43 = x42;
	assign y44 = x43;
	assign y45 = x44;
	assign y46 = x45;
	assign y47 = x46;
	assign y48 = x47;
	assign y49 = x48;
	assign y50 = x49;
	assign y51 = x50;
	assign y52 = x51;
	assign y53 = x52;
	assign y54 = x53;
	assign y55 = x54;
	assign y56 = x55;
	assign y57 = x56;
	assign y58 = x57;
	assign y59 = x58;
	assign y60 = x59;
	assign y61 = x60;
	assign y62 = x61;
	assign y63 = x62;
	assign y64 = x63;
	assign y65 = x64;
	assign y66 = x65;
	assign y67 = x66;
	assign y68 = x67;
	assign y69 = x68;
	assign y70 = x69;
	assign y71 = x70;
	assign y72 = x71;
	assign y73 = x72;
	assign y74 = x73;
	assign y75 = x74;
	assign y76 = x75;
	assign y77 = x76;
	assign y78 = x77;
	assign y79 = x78;
	assign y80 = x79;
	assign y81 = x80;
	assign y82 = x81;
	assign y83 = x82;
	assign y84 = x83;
	assign y85 = x84;
	assign y86 = x85;
	assign y87 = x86;
	assign y88 = x87;
	assign y89 = x88;
	assign y90 = x89;
	assign y91 = x90;
	assign y92 = x91;
	assign y93 = x92;
	assign y94 = x93;
	assign y95 = x94;
	assign y96 = x95;
	assign y97 = x96;
	assign y98 = x97;
	assign y99 = x98;
	assign y100 = x99;
	assign y101 = x100;
	assign y102 = x101;
	assign y103 = x102;
	assign y104 = x103;
	assign y105 = x104;
	assign y106 = x105;
	assign y107 = x106;
	assign y108 = x107;
	assign y109 = x108;
	assign y110 = x109;
	assign y111 = x110;
	assign y112 = x111;
	assign y113 = x112;
	assign y114 = x113;
	assign y115 = x114;
	assign y116 = x115;
	assign y117 = x116;
	assign y118 = x117;
	assign y119 = x118;
	assign y120 = x119;
	assign y121 = x120;
	assign y122 = x121;
	assign y123 = x122;
	assign y124 = x123;
	assign y125 = x124;
	assign y126 = x125;
	assign y127 = x126;
	assign y128 = x127;
	assign y129 = x128;
	assign y130 = x129;
	assign y131 = x130;
	assign y132 = x131;
	assign y133 = x132;
	assign y134 = x133;
	assign y135 = x134;
	assign y136 = x135;
	assign y137 = x136;
	assign y138 = x137;
	assign y139 = x138;
	assign y140 = x139;
	assign y141 = x140;
	assign y142 = x141;
	assign y143 = x142;
	assign y144 = x143;
	assign y145 = x144;
	assign y146 = x145;
	assign y147 = x146;
	assign y148 = x147;
	assign y149 = x148;
	assign y150 = x149;
	assign y151 = x150;
	assign y152 = x151;
	assign y153 = x152;
	assign y154 = x153;
	assign y155 = x154;
	assign y156 = x155;
	assign y157 = x156;
	assign y158 = x157;
	assign y159 = x158;
	assign y160 = x159;
	assign y161 = x160;
	assign y162 = x161;
	assign y163 = x162;
	assign y164 = x163;
	assign y165 = x164;
	assign y166 = x165;
	assign y167 = x166;
	assign y168 = x167;
	assign y169 = x168;
	assign y170 = x169;
	assign y171 = x170;
	assign y172 = x171;
	assign y173 = x172;
	assign y174 = x173;
	assign y175 = x174;
	assign y176 = x175;
	assign y177 = x176;
	assign y178 = x177;
	assign y179 = x178;
	assign y180 = x179;
	assign y181 = x180;
	assign y182 = x181;
	assign y183 = x182;
	assign y184 = x183;
	assign y185 = x184;
	assign y186 = x185;
	assign y187 = x186;
	assign y188 = x187;
	assign y189 = x188;
	assign y190 = x189;
	assign y191 = x190;
	assign y192 = x191;
	assign y193 = x192;
	assign y194 = x193;
	assign y195 = x194;
	assign y196 = x195;
	assign y197 = x196;
	assign y198 = x197;
	assign y199 = x198;
	assign y200 = x199;
	assign y201 = x200;
	assign y202 = x201;
	assign y203 = x202;
	assign y204 = x203;
	assign y205 = x204;
	assign y206 = x205;
	assign y207 = x206;
	assign y208 = x207;
	assign y209 = x208;
	assign y210 = x209;
	assign y211 = x210;
	assign y212 = x211;
	assign y213 = x212;
	assign y214 = x213;
	assign y215 = x214;
	assign y216 = x215;
	assign y217 = x216;
	assign y218 = x217;
	assign y219 = x218;
	assign y220 = x219;
	assign y221 = x220;
	assign y222 = x221;
	assign y223 = x222;
	assign y224 = x223;
	assign y225 = x224;
	assign y226 = x225;
	assign y227 = x226;
	assign y228 = x227;
	assign y229 = x228;
	assign y230 = x229;
	assign y231 = x230;
	assign y232 = x231;
	assign y233 = x232;
	assign y234 = x233;
	assign y235 = x234;
	assign y236 = x235;
	assign y237 = x236;
	assign y238 = x237;
	assign y239 = x238;
	assign y240 = x239;
	assign y241 = x240;
	assign y242 = x241;
	assign y243 = x242;
	assign y244 = x243;
	assign y245 = x244;
	assign y246 = x245;
	assign y247 = x246;
	assign y248 = x247;
	assign y249 = x248;
	assign y250 = x249;
	assign y251 = x250;
	assign y252 = x251;
	assign y253 = x252;
	assign y254 = x253;
	assign y255 = x254;
	assign y256 = x255;
	assign y257 = x256;
	assign y258 = x257;
	assign y259 = x258;
	assign y260 = x259;
	assign y261 = x260;
	assign y262 = x261;
	assign y263 = x262;
	assign y264 = x263;
	assign y265 = x264;
	assign y266 = x265;
	assign y267 = x266;
	assign y268 = x267;
	assign y269 = x268;
	assign y270 = x269;
	assign y271 = x270;
	assign y272 = x271;
	assign y273 = x272;
	assign y274 = x273;
	assign y275 = x274;
	assign y276 = x275;
	assign y277 = x276;
	assign y278 = x277;
	assign y279 = x278;
	assign y280 = x279;
	assign y281 = x280;
	assign y282 = x281;
	assign y283 = x282;
	assign y284 = x283;
	assign y285 = x284;
	assign y286 = x285;
	assign y287 = x286;
	assign y288 = x287;
	assign y289 = x288;
	assign y290 = x289;
	assign y291 = x290;
	assign y292 = x291;
	assign y293 = x292;
	assign y294 = x293;
	assign y295 = x294;
	assign y296 = x295;
	assign y297 = x296;
	assign y298 = x297;
	assign y299 = x298;
	assign y300 = x299;
	assign y301 = x300;
	assign y302 = x301;
	assign y303 = x302;
	assign y304 = x303;
	assign y305 = x304;
	assign y306 = x305;
	assign y307 = x306;
	assign y308 = x307;
	assign y309 = x308;
	assign y310 = x309;
	assign y311 = x310;
	assign y312 = x311;
	assign y313 = x312;
	assign y314 = x313;
	assign y315 = x314;
	assign y316 = x315;
	assign y317 = x316;
	assign y318 = x317;
	assign y319 = x318;
	assign y320 = x319;
	assign y321 = x320;
	assign y322 = x321;
	assign y323 = x322;
	assign y324 = x323;
	assign y325 = x324;
	assign y326 = x325;
	assign y327 = x326;
	assign y328 = x327;
	assign y329 = x328;
	assign y330 = x329;
	assign y331 = x330;
	assign y332 = x331;
	assign y333 = x332;
	assign y334 = x333;
	assign y335 = x334;
	assign y336 = x335;
	assign y337 = x336;
	assign y338 = x337;
	assign y339 = x338;
	assign y340 = x339;
	assign y341 = x340;
	assign y342 = x341;
	assign y343 = x342;
	assign y344 = x343;
	assign y345 = x344;
	assign y346 = x345;
	assign y347 = x346;
	assign y348 = x347;
	assign y349 = x348;
	assign y350 = x349;
	assign y351 = x350;
	assign y352 = x351;
	assign y353 = x352;
	assign y354 = x353;
	assign y355 = x354;
	assign y356 = x355;
	assign y357 = x356;
	assign y358 = x357;
	assign y359 = x358;
	assign y360 = x359;
	assign y361 = x360;
	assign y362 = x361;
	assign y363 = x362;
	assign y364 = x363;
	assign y365 = x364;
	assign y366 = x365;
	assign y367 = x366;
	assign y368 = x367;
	assign y369 = x368;
	assign y370 = x369;
	assign y371 = x370;
	assign y372 = x371;
	assign y373 = x372;
	assign y374 = x373;
	assign y375 = x374;
	assign y376 = x375;
	assign y377 = x376;
	assign y378 = x377;
	assign y379 = x378;
	assign y380 = x379;
	assign y381 = x380;
	assign y382 = x381;
	assign y383 = x382;
	assign y384 = x383;
	assign y385 = x384;
	assign y386 = x385;
	assign y387 = x386;
	assign y388 = x387;
	assign y389 = x388;
	assign y390 = x389;
	assign y391 = x390;
	assign y392 = x391;
	assign y393 = x392;
	assign y394 = x393;
	assign y395 = x394;
	assign y396 = x395;
	assign y397 = x396;
	assign y398 = x397;
	assign y399 = x398;
	assign y400 = x399;
	assign y401 = x400;
	assign y402 = x401;
	assign y403 = x402;
	assign y404 = x403;
	assign y405 = x404;
	assign y406 = x405;
	assign y407 = x406;
	assign y408 = x407;
	assign y409 = x408;
	assign y410 = x409;
	assign y411 = x410;
	assign y412 = x411;
	assign y413 = x412;
	assign y414 = x413;
	assign y415 = x414;
	assign y416 = x415;
	assign y417 = x416;
	assign y418 = x417;
	assign y419 = x418;
	assign y420 = x419;
	assign y421 = x420;
	assign y422 = x421;
	assign y423 = x422;
	assign y424 = x423;
	assign y425 = x424;
	assign y426 = x425;
	assign y427 = x426;
	assign y428 = x427;
	assign y429 = x428;
	assign y430 = x429;
	assign y431 = x430;
	assign y432 = x431;
	assign y433 = x432;
	assign y434 = x433;
	assign y435 = x434;
	assign y436 = x435;
	assign y437 = x436;
	assign y438 = x437;
	assign y439 = x438;
	assign y440 = x439;
	assign y441 = x440;
	assign y442 = x441;
	assign y443 = x442;
	assign y444 = x443;
	assign y445 = x444;
	assign y446 = x445;
	assign y447 = x446;
	always @(posedge clk)
		if (rst)
			d0 <= rst_val[0];
		else if (prog)
			d0 <= seed[0];
		else if (en)
			d0 <= x447;
	assign y0 = d0;
	assign x0a = y0;
	assign x21a = y0;
	assign x1a = y1;
	assign x22a = y1;
	assign x2a = y2;
	assign x23a = y2;
	assign x3a = y3;
	assign x24a = y3;
	assign x4a = y4;
	assign x25a = y4;
	assign x5a = y5;
	assign x26a = y5;
	assign x6a = y6;
	assign x27a = y6;
	assign x7a = y7;
	assign x28a = y7;
	assign x8a = y8;
	assign x29a = y8;
	assign x9a = y9;
	assign x30a = y9;
	assign x10a = y10;
	assign x31a = y10;
	assign x11a = y11;
	assign x32a = y11;
	assign x12a = y12;
	assign x33a = y12;
	assign x13a = y13;
	assign x34a = y13;
	assign x14a = y14;
	assign x35a = y14;
	assign x15a = y15;
	assign x36a = y15;
	assign x16a = y16;
	assign x37a = y16;
	assign x17a = y17;
	assign x38a = y17;
	assign x18a = y18;
	assign x39a = y18;
	assign x19a = y19;
	assign x40a = y19;
	assign x20a = y20;
	assign x41a = y20;
	assign x21b = y21;
	assign x42a = y21;
	assign x22b = y22;
	assign x43a = y22;
	assign x23b = y23;
	assign x44a = y23;
	assign x24b = y24;
	assign x45a = y24;
	assign x25b = y25;
	assign x46a = y25;
	assign x26b = y26;
	assign x47a = y26;
	assign x27b = y27;
	assign x48a = y27;
	assign x28b = y28;
	assign x49a = y28;
	assign x29b = y29;
	assign x50a = y29;
	assign x30b = y30;
	assign x51a = y30;
	assign x31b = y31;
	assign x52a = y31;
	assign x32b = y32;
	assign x53a = y32;
	assign x33b = y33;
	assign x54a = y33;
	assign x34b = y34;
	assign x55a = y34;
	assign x35b = y35;
	assign x56a = y35;
	assign x36b = y36;
	assign x57a = y36;
	assign x37b = y37;
	assign x58a = y37;
	assign x38b = y38;
	assign x59a = y38;
	assign x39b = y39;
	assign x60a = y39;
	assign x40b = y40;
	assign x61a = y40;
	assign x41b = y41;
	assign x62a = y41;
	assign x42b = y42;
	assign x63a = y42;
	assign x43b = y43;
	assign x64a = y43;
	assign x44b = y44;
	assign x65a = y44;
	assign x45b = y45;
	assign x66a = y45;
	assign x46b = y46;
	assign x67a = y46;
	assign x47b = y47;
	assign x68a = y47;
	assign x48b = y48;
	assign x69a = y48;
	assign x49b = y49;
	assign x70a = y49;
	assign x50b = y50;
	assign x71a = y50;
	assign x51b = y51;
	assign x72a = y51;
	assign x52b = y52;
	assign x73a = y52;
	assign x53b = y53;
	assign x74a = y53;
	assign x54b = y54;
	assign x75a = y54;
	assign x55b = y55;
	assign x76a = y55;
	assign x56b = y56;
	assign x77a = y56;
	assign x57b = y57;
	assign x78a = y57;
	assign x58b = y58;
	assign x79a = y58;
	assign x59b = y59;
	assign x80a = y59;
	assign x60b = y60;
	assign x81a = y60;
	assign x61b = y61;
	assign x82a = y61;
	assign x62b = y62;
	assign x83a = y62;
	assign x63b = y63;
	assign x84a = y63;
	assign x64b = y64;
	assign x85a = y64;
	assign x65b = y65;
	assign x86a = y65;
	assign x66b = y66;
	assign x87a = y66;
	assign x67b = y67;
	assign x88a = y67;
	assign x68b = y68;
	assign x89a = y68;
	assign x69b = y69;
	assign x90a = y69;
	assign x70b = y70;
	assign x91a = y70;
	assign x71b = y71;
	assign x92a = y71;
	assign x72b = y72;
	assign x93a = y72;
	assign x73b = y73;
	assign x94a = y73;
	assign x74b = y74;
	assign x95a = y74;
	assign x75b = y75;
	assign x96a = y75;
	assign x76b = y76;
	assign x97a = y76;
	assign x77b = y77;
	assign x98a = y77;
	assign x78b = y78;
	assign x99a = y78;
	assign x79b = y79;
	assign x100a = y79;
	assign x80b = y80;
	assign x101a = y80;
	assign x81b = y81;
	assign x102a = y81;
	assign x82b = y82;
	assign x103a = y82;
	assign x83b = y83;
	assign x104a = y83;
	assign x84b = y84;
	assign x105a = y84;
	assign x85b = y85;
	assign x106a = y85;
	assign x86b = y86;
	assign x107a = y86;
	assign x87b = y87;
	assign x108a = y87;
	assign x88b = y88;
	assign x109a = y88;
	assign x89b = y89;
	assign x110a = y89;
	assign x90b = y90;
	assign x111a = y90;
	assign x91b = y91;
	assign x112a = y91;
	assign x92b = y92;
	assign x113a = y92;
	assign x93b = y93;
	assign x114a = y93;
	assign x94b = y94;
	assign x115a = y94;
	assign x95b = y95;
	assign x116a = y95;
	assign x96b = y96;
	assign x117a = y96;
	assign x97b = y97;
	assign x118a = y97;
	assign x98b = y98;
	assign x119a = y98;
	assign x99b = y99;
	assign x120a = y99;
	assign x100b = y100;
	assign x121a = y100;
	assign x101b = y101;
	assign x122a = y101;
	assign x102b = y102;
	assign x123a = y102;
	assign x103b = y103;
	assign x124a = y103;
	assign x104b = y104;
	assign x125a = y104;
	assign x105b = y105;
	assign x126a = y105;
	assign x106b = y106;
	assign x127a = y106;
	assign x107b = y107;
	assign x128a = y107;
	assign x108b = y108;
	assign x129a = y108;
	assign x109b = y109;
	assign x130a = y109;
	assign x110b = y110;
	assign x131a = y110;
	assign x111b = y111;
	assign x132a = y111;
	assign x112b = y112;
	assign x133a = y112;
	assign x113b = y113;
	assign x134a = y113;
	assign x114b = y114;
	assign x135a = y114;
	assign x115b = y115;
	assign x136a = y115;
	assign x116b = y116;
	assign x137a = y116;
	assign x117b = y117;
	assign x138a = y117;
	assign x118b = y118;
	assign x139a = y118;
	assign x119b = y119;
	assign x140a = y119;
	assign x120b = y120;
	assign x141a = y120;
	assign x121b = y121;
	assign x142a = y121;
	assign x122b = y122;
	assign x143a = y122;
	assign x123b = y123;
	assign x144a = y123;
	assign x124b = y124;
	assign x145a = y124;
	assign x125b = y125;
	assign x146a = y125;
	assign x126b = y126;
	assign x147a = y126;
	assign x127b = y127;
	assign x148a = y127;
	assign x128b = y128;
	assign x149a = y128;
	assign x129b = y129;
	assign x150a = y129;
	assign x130b = y130;
	assign x151a = y130;
	assign x131b = y131;
	assign x152a = y131;
	assign x132b = y132;
	assign x153a = y132;
	assign x133b = y133;
	assign x154a = y133;
	assign x134b = y134;
	assign x155a = y134;
	assign x135b = y135;
	assign x156a = y135;
	assign x136b = y136;
	assign x157a = y136;
	assign x137b = y137;
	assign x158a = y137;
	assign x138b = y138;
	assign x159a = y138;
	assign x139b = y139;
	assign x160a = y139;
	assign x140b = y140;
	assign x161a = y140;
	assign x141b = y141;
	assign x162a = y141;
	assign x142b = y142;
	assign x163a = y142;
	assign x143b = y143;
	assign x164a = y143;
	assign x144b = y144;
	assign x165a = y144;
	assign x145b = y145;
	assign x166a = y145;
	assign x146b = y146;
	assign x167a = y146;
	assign x147b = y147;
	assign x168a = y147;
	assign x148b = y148;
	assign x169a = y148;
	assign x149b = y149;
	assign x170a = y149;
	assign x150b = y150;
	assign x171a = y150;
	assign x151b = y151;
	assign x172a = y151;
	assign x152b = y152;
	assign x173a = y152;
	assign x153b = y153;
	assign x174a = y153;
	assign x154b = y154;
	assign x175a = y154;
	assign x155b = y155;
	assign x176a = y155;
	assign x156b = y156;
	assign x177a = y156;
	assign x157b = y157;
	assign x178a = y157;
	assign x158b = y158;
	assign x179a = y158;
	assign x159b = y159;
	assign x180a = y159;
	assign x160b = y160;
	assign x181a = y160;
	assign x161b = y161;
	assign x182a = y161;
	assign x162b = y162;
	assign x183a = y162;
	assign x163b = y163;
	assign x184a = y163;
	assign x164b = y164;
	assign x185a = y164;
	assign x165b = y165;
	assign x186a = y165;
	assign x166b = y166;
	assign x187a = y166;
	assign x167b = y167;
	assign x188a = y167;
	assign x168b = y168;
	assign x189a = y168;
	assign x169b = y169;
	assign x190a = y169;
	assign x170b = y170;
	assign x191a = y170;
	assign x171b = y171;
	assign x192a = y171;
	assign x172b = y172;
	assign x193a = y172;
	assign x173b = y173;
	assign x194a = y173;
	assign x174b = y174;
	assign x195a = y174;
	assign x175b = y175;
	assign x196a = y175;
	assign x176b = y176;
	assign x197a = y176;
	assign x177b = y177;
	assign x198a = y177;
	assign x178b = y178;
	assign x199a = y178;
	assign x179b = y179;
	assign x200a = y179;
	assign x180b = y180;
	assign x201a = y180;
	assign x181b = y181;
	assign x202a = y181;
	assign x182b = y182;
	assign x203a = y182;
	assign x183b = y183;
	assign x204a = y183;
	assign x184b = y184;
	assign x205a = y184;
	assign x185b = y185;
	assign x206a = y185;
	assign x186b = y186;
	assign x207a = y186;
	assign x187b = y187;
	assign x208a = y187;
	assign x188b = y188;
	assign x209a = y188;
	assign x189b = y189;
	assign x210a = y189;
	assign x190b = y190;
	assign x211a = y190;
	assign x191b = y191;
	assign x212a = y191;
	assign x192b = y192;
	assign x213a = y192;
	assign x193b = y193;
	assign x214a = y193;
	assign x194b = y194;
	assign x215a = y194;
	assign x195b = y195;
	assign x216a = y195;
	assign x196b = y196;
	assign x217a = y196;
	assign x197b = y197;
	assign x218a = y197;
	assign x198b = y198;
	assign x219a = y198;
	assign x199b = y199;
	assign x220a = y199;
	assign x200b = y200;
	assign x221a = y200;
	assign x201b = y201;
	assign x222a = y201;
	assign x202b = y202;
	assign x223a = y202;
	assign x203b = y203;
	assign x224a = y203;
	assign x204b = y204;
	assign x225a = y204;
	assign x205b = y205;
	assign x226a = y205;
	assign x206b = y206;
	assign x227a = y206;
	assign x207b = y207;
	assign x228a = y207;
	assign x208b = y208;
	assign x229a = y208;
	assign x209b = y209;
	assign x230a = y209;
	assign x210b = y210;
	assign x231a = y210;
	assign x211b = y211;
	assign x232a = y211;
	assign x212b = y212;
	assign x233a = y212;
	assign x213b = y213;
	assign x234a = y213;
	assign x214b = y214;
	assign x235a = y214;
	assign x215b = y215;
	assign x236a = y215;
	assign x216b = y216;
	assign x237a = y216;
	assign x217b = y217;
	assign x238a = y217;
	assign x218b = y218;
	assign x239a = y218;
	assign x219b = y219;
	assign x240a = y219;
	assign x220b = y220;
	assign x241a = y220;
	assign x221b = y221;
	assign x242a = y221;
	assign x222b = y222;
	assign x243a = y222;
	assign x223b = y223;
	assign x244a = y223;
	assign x224b = y224;
	assign x245a = y224;
	assign x225b = y225;
	assign x246a = y225;
	assign x226b = y226;
	assign x247a = y226;
	assign x227b = y227;
	assign x248a = y227;
	assign x228b = y228;
	assign x249a = y228;
	assign x229b = y229;
	assign x250a = y229;
	assign x230b = y230;
	assign x251a = y230;
	assign x231b = y231;
	assign x252a = y231;
	assign x232b = y232;
	assign x253a = y232;
	assign x233b = y233;
	assign x254a = y233;
	assign x234b = y234;
	assign x255a = y234;
	assign x235b = y235;
	assign x256a = y235;
	assign x236b = y236;
	assign x257a = y236;
	assign x237b = y237;
	assign x258a = y237;
	assign x238b = y238;
	assign x259a = y238;
	assign x239b = y239;
	assign x260a = y239;
	assign x240b = y240;
	assign x261a = y240;
	assign x241b = y241;
	assign x262a = y241;
	assign x242b = y242;
	assign x263a = y242;
	assign x243b = y243;
	assign x264a = y243;
	assign x244b = y244;
	assign x265a = y244;
	assign x245b = y245;
	assign x266a = y245;
	assign x246b = y246;
	assign x267a = y246;
	assign x247b = y247;
	assign x268a = y247;
	assign x248b = y248;
	assign x269a = y248;
	assign x249b = y249;
	assign x270a = y249;
	assign x250b = y250;
	assign x271a = y250;
	assign x251b = y251;
	assign x272a = y251;
	assign x252b = y252;
	assign x273a = y252;
	assign x253b = y253;
	assign x274a = y253;
	assign x254b = y254;
	assign x275a = y254;
	assign x255b = y255;
	assign x276a = y255;
	assign x256b = y256;
	assign x277a = y256;
	assign x257b = y257;
	assign x278a = y257;
	assign x258b = y258;
	assign x279a = y258;
	assign x259b = y259;
	assign x280a = y259;
	assign x260b = y260;
	assign x281a = y260;
	assign x261b = y261;
	assign x282a = y261;
	assign x262b = y262;
	assign x283a = y262;
	assign x263b = y263;
	assign x284a = y263;
	assign x264b = y264;
	assign x285a = y264;
	assign x265b = y265;
	assign x286a = y265;
	assign x266b = y266;
	assign x287a = y266;
	assign x267b = y267;
	assign x288a = y267;
	assign x268b = y268;
	assign x289a = y268;
	assign x269b = y269;
	assign x290a = y269;
	assign x270b = y270;
	assign x291a = y270;
	assign x271b = y271;
	assign x292a = y271;
	assign x272b = y272;
	assign x293a = y272;
	assign x273b = y273;
	assign x294a = y273;
	assign x274b = y274;
	assign x295a = y274;
	assign x275b = y275;
	assign x296a = y275;
	assign x276b = y276;
	assign x297a = y276;
	assign x277b = y277;
	assign x298a = y277;
	assign x278b = y278;
	assign x299a = y278;
	assign x279b = y279;
	assign x300a = y279;
	assign x280b = y280;
	assign x301a = y280;
	assign x281b = y281;
	assign x302a = y281;
	assign x282b = y282;
	assign x303a = y282;
	assign x283b = y283;
	assign x304a = y283;
	assign x284b = y284;
	assign x305a = y284;
	assign x285b = y285;
	assign x306a = y285;
	assign x286b = y286;
	assign x307a = y286;
	assign x287b = y287;
	assign x308a = y287;
	assign x288b = y288;
	assign x309a = y288;
	assign x289b = y289;
	assign x310a = y289;
	assign x290b = y290;
	assign x311a = y290;
	assign x291b = y291;
	assign x312a = y291;
	assign x292b = y292;
	assign x313a = y292;
	assign x293b = y293;
	assign x314a = y293;
	assign x294b = y294;
	assign x315a = y294;
	assign x295b = y295;
	assign x316a = y295;
	assign x296b = y296;
	assign x317a = y296;
	assign x297b = y297;
	assign x318a = y297;
	assign x298b = y298;
	assign x319a = y298;
	assign x299b = y299;
	assign x320a = y299;
	assign x300b = y300;
	assign x321a = y300;
	assign x301b = y301;
	assign x322a = y301;
	assign x302b = y302;
	assign x323a = y302;
	assign x303b = y303;
	assign x324a = y303;
	assign x304b = y304;
	assign x325a = y304;
	assign x305b = y305;
	assign x326a = y305;
	assign x306b = y306;
	assign x327a = y306;
	assign x307b = y307;
	assign x328a = y307;
	assign x308b = y308;
	assign x329a = y308;
	assign x309b = y309;
	assign x330a = y309;
	assign x310b = y310;
	assign x331a = y310;
	assign x311b = y311;
	assign x332a = y311;
	assign x312b = y312;
	assign x333a = y312;
	assign x313b = y313;
	assign x334a = y313;
	assign x314b = y314;
	assign x335a = y314;
	assign x315b = y315;
	assign x336a = y315;
	assign x316b = y316;
	assign x337a = y316;
	assign x317b = y317;
	assign x338a = y317;
	assign x318b = y318;
	assign x339a = y318;
	assign x319b = y319;
	assign x340a = y319;
	assign x320b = y320;
	assign x341a = y320;
	assign x321b = y321;
	assign x342a = y321;
	assign x322b = y322;
	assign x343a = y322;
	assign x323b = y323;
	assign x344a = y323;
	assign x324b = y324;
	assign x345a = y324;
	assign x325b = y325;
	assign x346a = y325;
	assign x326b = y326;
	assign x347a = y326;
	assign x327b = y327;
	assign x348a = y327;
	assign x328b = y328;
	assign x349a = y328;
	assign x329b = y329;
	assign x350a = y329;
	assign x330b = y330;
	assign x351a = y330;
	assign x331b = y331;
	assign x352a = y331;
	assign x332b = y332;
	assign x353a = y332;
	assign x333b = y333;
	assign x354a = y333;
	assign x334b = y334;
	assign x355a = y334;
	assign x335b = y335;
	assign x356a = y335;
	assign x336b = y336;
	assign x357a = y336;
	assign x337b = y337;
	assign x358a = y337;
	assign x338b = y338;
	assign x359a = y338;
	assign x339b = y339;
	assign x360a = y339;
	assign x340b = y340;
	assign x361a = y340;
	assign x341b = y341;
	assign x362a = y341;
	assign x342b = y342;
	assign x363a = y342;
	assign x343b = y343;
	assign x364a = y343;
	assign x344b = y344;
	assign x365a = y344;
	assign x345b = y345;
	assign x366a = y345;
	assign x346b = y346;
	assign x367a = y346;
	assign x347b = y347;
	assign x368a = y347;
	assign x348b = y348;
	assign x369a = y348;
	assign x349b = y349;
	assign x370a = y349;
	assign x350b = y350;
	assign x371a = y350;
	assign x351b = y351;
	assign x372a = y351;
	assign x352b = y352;
	assign x373a = y352;
	assign x353b = y353;
	assign x374a = y353;
	assign x354b = y354;
	assign x375a = y354;
	assign x355b = y355;
	assign x376a = y355;
	assign x356b = y356;
	assign x377a = y356;
	assign x357b = y357;
	assign x378a = y357;
	assign x358b = y358;
	assign x379a = y358;
	assign x359b = y359;
	assign x380a = y359;
	assign x360b = y360;
	assign x381a = y360;
	assign x361b = y361;
	assign x382a = y361;
	assign x362b = y362;
	assign x383a = y362;
	assign x363b = y363;
	assign x384a = y363;
	assign x364b = y364;
	assign x385a = y364;
	assign x365b = y365;
	assign x386a = y365;
	assign x366b = y366;
	assign x387a = y366;
	assign x367b = y367;
	assign x388a = y367;
	assign x368b = y368;
	assign x389a = y368;
	assign x369b = y369;
	assign x390a = y369;
	assign x370b = y370;
	assign x391a = y370;
	assign x371b = y371;
	assign x392a = y371;
	assign x372b = y372;
	assign x393a = y372;
	assign x373b = y373;
	assign x394a = y373;
	assign x374b = y374;
	assign x395a = y374;
	assign x375b = y375;
	assign x396a = y375;
	assign x376b = y376;
	assign x397a = y376;
	assign x377b = y377;
	assign x398a = y377;
	assign x378b = y378;
	assign x399a = y378;
	assign x379b = y379;
	assign x400a = y379;
	assign x380b = y380;
	assign x401a = y380;
	assign x381b = y381;
	assign x402a = y381;
	assign x382b = y382;
	assign x403a = y382;
	assign x383b = y383;
	assign x404a = y383;
	assign x384b = y384;
	assign x405a = y384;
	assign x385b = y385;
	assign x406a = y385;
	assign x386b = y386;
	assign x407a = y386;
	assign x387b = y387;
	assign x408a = y387;
	assign x388b = y388;
	assign x409a = y388;
	assign x389b = y389;
	assign x410a = y389;
	assign x390b = y390;
	assign x411a = y390;
	assign x391b = y391;
	assign x412a = y391;
	assign x392b = y392;
	assign x413a = y392;
	assign x393b = y393;
	assign x414a = y393;
	assign x394b = y394;
	assign x415a = y394;
	assign x395b = y395;
	assign x416a = y395;
	assign x396b = y396;
	assign x417a = y396;
	assign x397b = y397;
	assign x418a = y397;
	assign x398b = y398;
	assign x419a = y398;
	assign x399b = y399;
	assign x420a = y399;
	assign x400b = y400;
	assign x421a = y400;
	assign x401b = y401;
	assign x422a = y401;
	assign x402b = y402;
	assign x423a = y402;
	assign x403b = y403;
	assign x424a = y403;
	assign x404b = y404;
	assign x425a = y404;
	assign x405b = y405;
	assign x426a = y405;
	assign x406b = y406;
	assign x427a = y406;
	assign x407b = y407;
	assign x428a = y407;
	assign x408b = y408;
	assign x429a = y408;
	assign x409b = y409;
	assign x430a = y409;
	assign x410b = y410;
	assign x431a = y410;
	assign x411b = y411;
	assign x432a = y411;
	assign x412b = y412;
	assign x433a = y412;
	assign x413b = y413;
	assign x434a = y413;
	assign x414b = y414;
	assign x435a = y414;
	assign x415b = y415;
	assign x436a = y415;
	assign x416b = y416;
	assign x437a = y416;
	assign x417b = y417;
	assign x438a = y417;
	assign x418b = y418;
	assign x439a = y418;
	assign x419b = y419;
	assign x440a = y419;
	assign x420b = y420;
	assign x441a = y420;
	assign x421b = y421;
	assign x442a = y421;
	assign x422b = y422;
	assign x443a = y422;
	assign x423b = y423;
	assign x444a = y423;
	assign x424b = y424;
	assign x445a = y424;
	assign x425b = y425;
	assign x446a = y425;
	assign x426b = y426;
	assign x447a = y426;
	assign x427b = y427;
	always @(posedge clk)
		if (rst)
			d1 <= rst_val[1];
		else if (prog)
			d1 <= seed[1];
		else if (en)
			d1 <= y427;
	assign x0b = d1;
	assign x428b = y428;
	always @(posedge clk)
		if (rst)
			d2 <= rst_val[2];
		else if (prog)
			d2 <= seed[2];
		else if (en)
			d2 <= y428;
	assign x1b = d2;
	assign x429b = y429;
	always @(posedge clk)
		if (rst)
			d3 <= rst_val[3];
		else if (prog)
			d3 <= seed[3];
		else if (en)
			d3 <= y429;
	assign x2b = d3;
	assign x430b = y430;
	always @(posedge clk)
		if (rst)
			d4 <= rst_val[4];
		else if (prog)
			d4 <= seed[4];
		else if (en)
			d4 <= y430;
	assign x3b = d4;
	assign x431b = y431;
	always @(posedge clk)
		if (rst)
			d5 <= rst_val[5];
		else if (prog)
			d5 <= seed[5];
		else if (en)
			d5 <= y431;
	assign x4b = d5;
	assign x432b = y432;
	always @(posedge clk)
		if (rst)
			d6 <= rst_val[6];
		else if (prog)
			d6 <= seed[6];
		else if (en)
			d6 <= y432;
	assign x5b = d6;
	assign x433b = y433;
	always @(posedge clk)
		if (rst)
			d7 <= rst_val[7];
		else if (prog)
			d7 <= seed[7];
		else if (en)
			d7 <= y433;
	assign x6b = d7;
	assign x434b = y434;
	always @(posedge clk)
		if (rst)
			d8 <= rst_val[8];
		else if (prog)
			d8 <= seed[8];
		else if (en)
			d8 <= y434;
	assign x7b = d8;
	assign x435b = y435;
	always @(posedge clk)
		if (rst)
			d9 <= rst_val[9];
		else if (prog)
			d9 <= seed[9];
		else if (en)
			d9 <= y435;
	assign x8b = d9;
	assign x436b = y436;
	always @(posedge clk)
		if (rst)
			d10 <= rst_val[10];
		else if (prog)
			d10 <= seed[10];
		else if (en)
			d10 <= y436;
	assign x9b = d10;
	assign x437b = y437;
	always @(posedge clk)
		if (rst)
			d11 <= rst_val[11];
		else if (prog)
			d11 <= seed[11];
		else if (en)
			d11 <= y437;
	assign x10b = d11;
	assign x438b = y438;
	always @(posedge clk)
		if (rst)
			d12 <= rst_val[12];
		else if (prog)
			d12 <= seed[12];
		else if (en)
			d12 <= y438;
	assign x11b = d12;
	assign x439b = y439;
	always @(posedge clk)
		if (rst)
			d13 <= rst_val[13];
		else if (prog)
			d13 <= seed[13];
		else if (en)
			d13 <= y439;
	assign x12b = d13;
	assign x440b = y440;
	always @(posedge clk)
		if (rst)
			d14 <= rst_val[14];
		else if (prog)
			d14 <= seed[14];
		else if (en)
			d14 <= y440;
	assign x13b = d14;
	assign x441b = y441;
	always @(posedge clk)
		if (rst)
			d15 <= rst_val[15];
		else if (prog)
			d15 <= seed[15];
		else if (en)
			d15 <= y441;
	assign x14b = d15;
	assign x442b = y442;
	always @(posedge clk)
		if (rst)
			d16 <= rst_val[16];
		else if (prog)
			d16 <= seed[16];
		else if (en)
			d16 <= y442;
	assign x15b = d16;
	assign x443b = y443;
	always @(posedge clk)
		if (rst)
			d17 <= rst_val[17];
		else if (prog)
			d17 <= seed[17];
		else if (en)
			d17 <= y443;
	assign x16b = d17;
	assign x444b = y444;
	always @(posedge clk)
		if (rst)
			d18 <= rst_val[18];
		else if (prog)
			d18 <= seed[18];
		else if (en)
			d18 <= y444;
	assign x17b = d18;
	assign x445b = y445;
	always @(posedge clk)
		if (rst)
			d19 <= rst_val[19];
		else if (prog)
			d19 <= seed[19];
		else if (en)
			d19 <= y445;
	assign x18b = d19;
	assign x446b = y446;
	always @(posedge clk)
		if (rst)
			d20 <= rst_val[20];
		else if (prog)
			d20 <= seed[20];
		else if (en)
			d20 <= y446;
	assign x19b = d20;
	assign x447b = y447;
	always @(posedge clk)
		if (rst)
			d21 <= rst_val[21];
		else if (prog)
			d21 <= seed[21];
		else if (en)
			d21 <= y447;
	assign x20b = d21;

	// Output assignment
	assign out = {y447,y446,y445,y444,y443,y442,y441,y440,y439,y438,y437,y436,y435,y434,y433,y432,y431,y430,y429,y428,y427,y426,y425,y424,y423,y422,y421,y420,y419,y418,y417,y416,y415,y414,y413,y412,y411,y410,y409,y408,y407,y406,y405,y404,y403,y402,y401,y400,y399,y398,y397,y396,y395,y394,y393,y392,y391,y390,y389,y388,y387,y386,y385,y384,y383,y382,y381,y380,y379,y378,y377,y376,y375,y374,y373,y372,y371,y370,y369,y368,y367,y366,y365,y364,y363,y362,y361,y360,y359,y358,y357,y356,y355,y354,y353,y352,y351,y350,y349,y348,y347,y346,y345,y344,y343,y342,y341,y340,y339,y338,y337,y336,y335,y334,y333,y332,y331,y330,y329,y328,y327,y326,y325,y324,y323,y322,y321,y320,y319,y318,y317,y316,y315,y314,y313,y312,y311,y310,y309,y308,y307,y306,y305,y304,y303,y302,y301,y300,y299,y298,y297,y296,y295,y294,y293,y292,y291,y290,y289,y288,y287,y286,y285,y284,y283,y282,y281,y280,y279,y278,y277,y276,y275,y274,y273,y272,y271,y270,y269,y268,y267,y266,y265,y264,y263,y262,y261,y260,y259,y258,y257,y256,y255,y254,y253,y252,y251,y250,y249,y248,y247,y246,y245,y244,y243,y242,y241,y240,y239,y238,y237,y236,y235,y234,y233,y232,y231,y230,y229,y228,y227,y226,y225,y224,y223,y222,y221,y220,y219,y218,y217,y216,y215,y214,y213,y212,y211,y210,y209,y208,y207,y206,y205,y204,y203,y202,y201,y200,y199,y198,y197,y196,y195,y194,y193,y192,y191,y190,y189,y188,y187,y186,y185,y184,y183,y182,y181,y180,y179,y178,y177,y176,y175,y174,y173,y172,y171,y170,y169,y168,y167,y166,y165,y164,y163,y162,y161,y160,y159,y158,y157,y156,y155,y154,y153,y152,y151,y150,y149,y148,y147,y146,y145,y144,y143,y142,y141,y140,y139,y138,y137,y136,y135,y134,y133,y132,y131,y130,y129,y128,y127,y126,y125,y124,y123,y122,y121,y120,y119,y118,y117,y116,y115,y114,y113,y112,y111,y110,y109,y108,y107,y106,y105,y104,y103,y102,y101,y100,y99,y98,y97,y96,y95,y94,y93,y92,y91,y90,y89,y88,y87,y86,y85,y84,y83,y82,y81,y80,y79,y78,y77,y76,y75,y74,y73,y72,y71,y70,y69,y68,y67,y66,y65,y64,y63,y62,y61,y60,y59,y58,y57,y56,y55,y54,y53,y52,y51,y50,y49,y48,y47,y46,y45,y44,y43,y42,y41,y40,y39,y38,y37,y36,y35,y34,y33,y32,y31,y30,y29,y28,y27,y26,y25,y24,y23,y22,y21,y20,y19,y18,y17,y16,y15,y14,y13,y12,y11,y10,y9,y8,y7,y6,y5,y4,y3,y2,y1,y0};

endmodule
